`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Lillia
// 
// Create Date: 2026/01/14 18:41:28
// Design Name: SD��ģ�ͣ�SPIЭ�飩
// Module Name: sd_model
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sd_model(
    input   wire    sd_clk,     // ����FPGA��SPIʱ��
    input   wire    sd_mosi,    // ����FPGA����������
    input   wire    sd_cs_n,    // ����FPGA��Ƭѡ�źţ�����Ч��
    output  reg     sd_miso     // ����FPGA���������
);

    // �洢���������
    // 169���� * 4096���� * 2�ֽ� = 1,384,448 �ֽڣ�һ��16λ������ռ�����ֽڣ�
    parameter   MEM_SIZE = 1384448; 
    reg [7:0]   mem[MEM_SIZE-1:0];  // 1byte == 8bits
 
    reg [47:0]  cmd_buffer;   
    reg [1:0]   STATE; 
    reg         is_acmd_prefix;     // ���ڱ�־��һ������ΪACMD  
    reg         stop_flag;          // ����ֹͣ������ȡ�ı�־λ
    reg [5:0]   rx_bit_cnt;         // ר�����ڽ�������ļ�����
    reg         start_multi_read;   // ���ڴ��������߼�
    reg         busy;               // ���ڱ�־�������ڽ���
    
    reg [5:0]   saved_idx;          // �����ݴ�ָ����
    reg [31:0]  saved_arg;          // �����ݴ��ַ����
    
    // ״̬����
    localparam  IDLE  = 2'b00,    // ���� 
                INIT  = 2'b01,    // ��ʼ��ʼ��
                READY = 2'b10;    // ��ʼ�������
                
    // ��ʼ����
    initial begin
        $readmemh("data_5band.txt", mem);
        sd_miso         = 1'b1;      
        STATE           = IDLE;
        is_acmd_prefix  = 0;
    end
    
    // ר�ŵĽ��ս��̣�ʼ�����У����ܷ��������Ӱ��
    always @(posedge sd_clk) begin
        if (sd_cs_n) begin     // ƬѡΪ1ʱΪ����
            rx_bit_cnt <= 0;
            cmd_buffer <= 48'b0;
            stop_flag <= 1'b0;
            start_multi_read <= 1'b0;
            busy <= 1'd0;
            
            saved_idx <= 6'd0;
            saved_arg <= 32'd0;
            // ��Ƭѡ���ߣ�ǿ����ֹ��������ȷ����λ
            disable send_data_sector;
            disable send_multi_data_blocks;
            disable send_r1;
        end else begin    // ƬѡΪ0ʱ������ʼ���
            if(!busy)
                if (rx_bit_cnt < 48) begin    // ����ʱ���߼�����������n��ʱ˵���Ѷ�ȡ��n��λ
                    cmd_buffer <= {cmd_buffer[46:0], sd_mosi};
                    rx_bit_cnt <= rx_bit_cnt + 1;
                end else begin    // ��ȡ�����һλ
                    rx_bit_cnt <= 0;
                    busy <= 1'd1;    // ��־����ʼ��֮���ܿ�ʼ����������cs���ߣ����·�������
                    handle_command(cmd_buffer);    // �����߼�״̬
                end
        end
    end
    
    // �������
    // ���ｫ����Ͳ�����Ϊȫ�֣��Ա㷢�Ͷ������ʱ���Ե���
    task handle_command(input [47:0] cmd);
        begin
            saved_idx = cmd[45:40];
            saved_arg = cmd[39:8];    // ��ȡ��������ΪSPI���ù�CRCУ�飬����Ͳ����ˣ�
            case(saved_idx)
                6'd0: begin
                    STATE = INIT;    // ����ΪCMD0ʱ˵����ʼ��ʼ��
                    send_r1(8'h01); 
                end
                
                6'd8: begin 
                    send_r7(8'h01, 32'h000001AA);
                end
                
                6'd55: begin 
                    is_acmd_prefix = 1;    // ���ߣ�˵����һ������������Ӧ������
                    send_r1(8'h01);
                end
                
                6'd41: begin 
                    if(is_acmd_prefix) begin    // ֻ������Ϊ����Ӧ���������Ӧ��������0x04
                        STATE = READY;    // ����Ϊ41ʱ˵����ʼ�����
                        send_r1(8'h00);   
                        is_acmd_prefix = 0;    // �����������״̬
                    end else 
                        send_r1(8'h04);
                end
                
                6'd17: begin 
                    if(STATE == READY)    // ��ʼ�����
                        send_data_sector(saved_arg);
                    else 
                        send_r1(8'h01);
                end
                
                6'd18: begin
                    if(STATE == READY) begin    // ��ʼ�����
                        stop_flag = 0;
                        saved_arg <= cmd[39:8];
                        start_multi_read = 1;    // ���������߼��������ﲻҪֱ�ӵ���    
                    end else
                        send_r1(8'h01);
                end
                
                6'd12: begin
                    stop_flag = 1; // �յ�ָֹͣ��޸ı�־λ����send_multi_data_blocks�˳�ѭ��
                end
                
                default: 
                    send_r1(8'h00);
            endcase
        end
    endtask
    
    // ���÷�������飬����Ӱ��cmd��ȡ
    always @(posedge sd_clk) begin
        if (start_multi_read) begin
            start_multi_read <= 0;
            send_multi_data_blocks(saved_arg); // ���÷�������
        end
    end
    
    // ��������
    task send_r1(input [7:0] r1_val);
        integer i;
        reg [7:0] temp_r1; // �����м��������Ϊ���벻��λ����
        begin
            temp_r1 = r1_val; 
            repeat(8) @(negedge sd_clk);    // �ֶ��ȴ�8��ʱ���½��أ�NCR�ӳ٣�ģ����ʵSD���Ĵ���ʱ�䣩
            for (i=0; i<8; i=i+1) begin
                sd_miso = temp_r1[7-i];
                @(negedge sd_clk);
                /* ��������һ��֮�����˼��
                   ִ������һ�β�����ȵ���һ��sd_clk���½����������߻�ѭ��
                   ʵ���Ͼ������½��ص�ʱ��׼������ȷ��miso�������ȶ�����
                   */
            end
            sd_miso = 1'b1;    // ���ݷ�����Ϻ���1
        end
    endtask

    task send_r7(input [7:0] r1_val, input [31:0] r7_val);
        integer i;
        reg [31:0] temp_r7;
        begin
            send_r1(r1_val);
            temp_r7 = r7_val;    // ������ֵ��miso��1��Ч����һ��ʱ���½����������32λ����
            for (i=31; i>=0; i=i-1) begin
                sd_miso = temp_r7[i];
                @(negedge sd_clk);
            end
            sd_miso = 1'b1;    // ���ݷ�����Ϻ���1
        end
    endtask
    
    // ���͵�������
    task send_data_sector(input [31:0] address);
        integer i, j;
        reg [7:0] target_byte;
        reg [31:0] real_byte_addr;
        reg [7:0] token; // �����м������� 0xFE
        begin
            send_r1(8'h00);
            repeat(16) @(negedge sd_clk);    // �ֶ��ȴ�16��ʱ���½��أ�NCR�ӳ٣�ģ����ʵSD����Ѱַʱ�䣩
            
            token = 8'hFE;    // ׼������ͷ��־
            for (i=7; i>=0; i=i-1) begin
                sd_miso = token[i];    // ��������ͷ
                @(negedge sd_clk);
            end

            real_byte_addr = address * 512;    // �������׸����ݵĵ�ַ
            for (i=0; i<512; i=i+1) begin
                if (real_byte_addr + i < MEM_SIZE)
                    target_byte = mem[real_byte_addr + i];    // ����Խ�����
                else
                    target_byte = 8'h00;

                for (j=7; j>=0; j=j-1) begin
                    sd_miso = target_byte[j];    // ѭ�������ֽڣ��ߵ��ͣ�
                    @(negedge sd_clk);
                end
            end

            repeat(16) begin
                sd_miso = 1'b1;    // ģ�ⷢ��CRCУ��ֵ0xFF��SPI�������Զ�����
                @(negedge sd_clk);
            end
        end
    endtask

    // ������������ ---
    task send_multi_data_blocks(input [31:0] start_address);
        integer i, j;
        reg [31:0] current_sector;
        reg [31:0] real_byte_addr;
        reg [7:0] target_byte;
        reg [7:0] token; // �����м������� 0xFE
        begin
            send_r1(8'h00); // ���� CMD18 ����Ӧ
            current_sector = start_address;
            
            // ֻҪû���յ�ֹͣ�źţ���һֱ����
            while (!stop_flag) begin
                // ���CS����ֹ��ѭ��
                if (sd_cs_n) begin
                     stop_flag = 1; 
                end
                repeat(8) @(negedge sd_clk); // ����ӳ�
                
                // 1. ������ʼ���� 0xFE
                token = 8'hFE;    // ׼������ͷ��־
                for (i=7; i>=0; i=i-1) begin
                    sd_miso = token[i];
                    @(negedge sd_clk);
                end

                // 2. ���� 512 �ֽ�����
                real_byte_addr = current_sector * 512;
                for (i=0; i<512; i=i+1) begin
                    if (real_byte_addr + i < MEM_SIZE)
                        target_byte = mem[real_byte_addr + i];
                    else
                        target_byte = 8'h00;

                    for (j=7; j>=0; j=j-1) begin
                        sd_miso = target_byte[j];
                        @(negedge sd_clk);
                    end
                end

                // 3. ���� 16 λ CRC (0xFFFF)
                repeat(16) begin
                    sd_miso = 1'b1;
                    @(negedge sd_clk);
                end
                
                // 4. ָ����һ������
                current_sector = current_sector + 1;
                
                // ���ؼ��߼������ڿ鷢����Ϻ󣬼���Ƿ��յ� CMD12
                // ����ڷ����ڼ� stop_flag �� handle_command �޸��ˣ�ѭ���ͻ��˳�
                // ע�⣺��ʵ�ʷ����У�����Task�������ģ���Ҫ��⵽CMD12��
                // ����FPGA�������������ݿ�֮��Ŀ����ڷ���ָ�
                if (current_sector * 512 >= MEM_SIZE) stop_flag = 1;
            end
            
            sd_miso = 1'b1; 
        end
    endtask
    
endmodule





