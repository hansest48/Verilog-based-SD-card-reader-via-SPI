`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Lillia
// 
// Create Date: 2026/01/15 17:51:34
// Design Name: ��ȡSD��������������
// Module Name: sd_read
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sd_read(
    input   wire    sd_clk,
    /* ����ʱ�ӣ������ն˲���
       ����SD�����ź�ʱ��ƫ�� */
    input   wire    sd_clk_i,
    input   wire    sd_rst_n,
    input   wire    sdinit_ok,  // ��ʼ���ɹ���־
    input   wire            addr_TVALID,  // ��ַ��Чλ
    input   wire    [31:0]  addr,         // ������ַ 
    
    input   wire    sd_miso,    // ����SD������������
    output  reg     sd_cs_n,    // ����SD����Ƭѡ�źţ�����Ч��
    output  reg     sd_mosi,    // ����SD�����������  
    
    output  reg         SectorData_TVALID,
    output  reg [15:0]  SectorData_TDATA,
    output  reg         SectorData_TLAST
    );
    
    // ״̬����
    localparam  IDLE        = 3'b000,    // ����
                WAIT_INIT   = 3'b001,    // �ȴ���ʼ��
                SEND_CMD    = 3'b010,    // ����48λ����
                WAIT_R1     = 3'b011,    // �ȴ�R1��Ӧ
                WAIT_TOKEN  = 3'b100,    // �ȴ���������0xFE
                READ_DATA   = 3'b101,    // ��ȡ512�ֽ�����
                READ_CRC    = 3'b110,    // ��ȡ16λCRC
                DONE        = 3'b111;    // ���ݽ������
                
    // SD��ָ�
    reg [47:0] CMD17;
    
    reg [2:0]  STATE;
    reg [5:0]  wait_cnt;    // ����ǰ�ȴ�
    reg        cmd_start;   // ���ʼλ
    reg [5:0]  bit_cnt;     // λ������
    reg [47:0] cmd_reg;     // ����Ĵ���
    reg [7:0]  res_reg;     // ��Ӧ���ռĴ���
    reg        receiving;   // ��Ӧ�����б�־λ       
    reg [8:0]  byte_cnt;    // 512�ֽڼ�����
    reg [7:0]  byte_data;   // �ֽ���װ�Ĵ���
    reg [7:0]  high_byte;   // 16λ���ݵĸ��ֽ��ݴ�
    reg        byte_sel;    // �ֽ�ѡ��1:���ֽ�, 0:���ֽڣ�������ƿ���������Ĵ������һ���ʺ���������ķ�����
    
    // ����ʱ�Ӳ���MISO������̬
    reg miso_d1;
    always @(posedge sd_clk_i) begin
        miso_d1 <= sd_miso;
    end
    
    // ״̬��
    always @(posedge sd_clk or negedge sd_rst_n) begin
        if (!sd_rst_n) begin
            STATE    <= IDLE;
            CMD17    <= 48'd0;
            wait_cnt <= 6'd0;
            cmd_start <= 1'd0;
            bit_cnt  <= 6'd0;
            cmd_reg  <= 48'd0;
            res_reg  <= 40'd0;
            receiving <= 'd0;
            
            sd_cs_n  <= 1'b1;
            sd_mosi  <= 1'b1;
            
            SectorData_TVALID <= 1'b0;
            SectorData_TDATA <= 16'b0;
            SectorData_TLAST <= 1'b0;
            
            byte_cnt  <= 9'd0;
            byte_data <= 8'd0;
            high_byte <= 8'd0;
            byte_sel  <= 1'b1;
            
        end else begin
            case(STATE)
                IDLE: begin
                    sd_cs_n <= 1'b1;    // ƬѡΪ1ʱΪ����
                    sd_mosi <= 1'b1;
                    SectorData_TVALID <= 1'b0;
                    SectorData_TLAST <= 1'b0;
                    STATE <= WAIT_INIT;
                end
                
                // 1 �ȴ���ʼ�����
                WAIT_INIT:
                    if(sdinit_ok)
                        STATE <= SEND_CMD;
                        
                // 2 �������48 bits��
                SEND_CMD: begin
                    if(addr_TVALID) begin
                        CMD17 <= {8'h51, addr, 8'hFF}; 
                        cmd_start <= 1'd1;
                    end
    
                    // ��������
                    if(cmd_start)
                        if (bit_cnt == 6'd0) begin
                            sd_cs_n <= 1'b0;    // ����Ƭѡ����ͬ����������
                            cmd_reg <= CMD17;
                            sd_mosi <= 0;
                            bit_cnt <= bit_cnt + 1'b1;
                        end else if(bit_cnt >= 1 && bit_cnt < 6'd48) begin    // ����48�������Զ�ת״̬����������������
                            sd_mosi <= cmd_reg[46];    // ѭ�������2λ����Ϊ��1λһ����0��ֻ��bit_cnt��1����ѭ����
                            cmd_reg <= {cmd_reg[46:0], 1'b1};
                            bit_cnt <= bit_cnt + 1'b1;
                        end else begin
                            cmd_start <= 1'd0;
                            bit_cnt <= 6'd0;
                            sd_mosi <= 1'b1;    // ������ͷ�mosi
                            STATE <= WAIT_R1; // ����ȴ���Ӧ״̬
                        end
                end
                
                // 3 �ȴ���Ӧ
                WAIT_R1: begin
                    if (miso_d1 == 1'b0 || receiving) begin
                        receiving <= 1'b1;
                        if (bit_cnt < 6'd8) begin
                            bit_cnt <= bit_cnt + 1'b1;
                            res_reg <= {res_reg[6:0], miso_d1};
                        end else begin
                            bit_cnt <= 6'd0;
                            receiving <= 1'b0;
                            if (res_reg == 8'h00)
                                STATE <= WAIT_TOKEN;    // �յ�R1����ʼ����������
                            else
                                STATE <= SEND_CMD;    // δ�յ�R1�����·���CMD
                        end
                    end
                end
                
                // 4 �ȴ�����ͷTOKEN��SD���м��һֱ����FF����⵽FE���һλ��0�Ϳ��Լ�����
                WAIT_TOKEN: begin
                    if (miso_d1 == 1'b0) begin // 0xFE�����һλ��0
                        STATE <= READ_DATA;
                        bit_cnt <= 6'd0;
                        byte_cnt <= 9'd0;
                        byte_sel <= 1'b1;
                    end
                end
                
                // 5 ��ȡ512�ֽڲ�תΪ16λ���
                READ_DATA: begin
                    if (bit_cnt < 6'd7) begin    // �ȶ�7λ�����һλ����ʱ��˳�㸳ֵ���ߵ�λ
                        byte_data <= {byte_data[6:0], miso_d1};
                        bit_cnt <= bit_cnt + 1'b1;
                    end else begin
                        bit_cnt <= 6'd0;
                        // �ֽڽ�����ɣ��ж��Ǹ�λ���ǵ�λ
                        if (byte_sel == 1'b1) begin
                            high_byte <= {byte_data[6:0], miso_d1};    // ����Ǹ�λ�ʹ�����
                            byte_sel <= 1'b0;
                        end else begin
                            SectorData_TDATA <= {high_byte, byte_data[6:0], miso_d1};    // ����ǵ�λ�ͺ͸�λ��ϲ����
                            SectorData_TVALID <= 1'b1;
                            byte_sel <= 1'b1;
                            if (byte_cnt == 511) 
                                SectorData_TLAST <= 1'b1;
                        end

                        if (byte_cnt < 511)
                            byte_cnt <= byte_cnt + 1'b1;    // �ڶ�ÿ���ֽ����һλʱ����
                        else begin
                            byte_cnt <= 9'd0;
                            STATE <= READ_CRC;
                        end
                    end
                end

                // 6 ��ȡ16λCRC������
                READ_CRC: begin
                    SectorData_TVALID <= 1'b0;
                    SectorData_TLAST <= 1'b0;
                    if (bit_cnt < 6'd15) begin
                        bit_cnt <= bit_cnt + 1'b1;
                    end else begin
                        bit_cnt <= 6'd0;
                        STATE <= DONE;
                    end
                end
                
                DONE: begin
                    sd_cs_n <= 1'b1;
                    STATE <= IDLE;
                end

                default: STATE <= IDLE;
            endcase   
        end 
    end       
endmodule



